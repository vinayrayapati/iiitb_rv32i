VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO iiitb_rv32i
  CLASS BLOCK ;
  FOREIGN iiitb_rv32i ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 650.000 ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END RN
  PIN WB_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 646.000 203.230 650.000 ;
    END
  END WB_OUT[0]
  PIN WB_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END WB_OUT[10]
  PIN WB_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 646.000 573.530 650.000 ;
    END
  END WB_OUT[11]
  PIN WB_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 646.000 55.110 650.000 ;
    END
  END WB_OUT[12]
  PIN WB_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 646.000 499.470 650.000 ;
    END
  END WB_OUT[13]
  PIN WB_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END WB_OUT[14]
  PIN WB_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END WB_OUT[15]
  PIN WB_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 411.440 650.000 412.040 ;
    END
  END WB_OUT[1]
  PIN WB_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END WB_OUT[2]
  PIN WB_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END WB_OUT[3]
  PIN WB_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 489.640 650.000 490.240 ;
    END
  END WB_OUT[4]
  PIN WB_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 333.240 650.000 333.840 ;
    END
  END WB_OUT[5]
  PIN WB_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END WB_OUT[6]
  PIN WB_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 646.000 425.410 650.000 ;
    END
  END WB_OUT[7]
  PIN WB_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 646.000 129.170 650.000 ;
    END
  END WB_OUT[8]
  PIN WB_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END WB_OUT[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 98.640 650.000 99.240 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 646.000 647.590 650.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 20.440 650.000 21.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 176.840 650.000 177.440 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 567.840 650.000 568.440 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 646.000 277.290 650.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 646.000 351.350 650.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 255.040 650.000 255.640 ;
    END
  END io_oeb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 636.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 636.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 636.565 ;
      LAYER met1 ;
        RECT 0.070 10.640 647.610 642.560 ;
      LAYER met2 ;
        RECT 0.100 645.720 54.550 646.000 ;
        RECT 55.390 645.720 128.610 646.000 ;
        RECT 129.450 645.720 202.670 646.000 ;
        RECT 203.510 645.720 276.730 646.000 ;
        RECT 277.570 645.720 350.790 646.000 ;
        RECT 351.630 645.720 424.850 646.000 ;
        RECT 425.690 645.720 498.910 646.000 ;
        RECT 499.750 645.720 572.970 646.000 ;
        RECT 573.810 645.720 647.030 646.000 ;
        RECT 0.100 4.280 647.580 645.720 ;
        RECT 0.650 4.000 73.870 4.280 ;
        RECT 74.710 4.000 147.930 4.280 ;
        RECT 148.770 4.000 221.990 4.280 ;
        RECT 222.830 4.000 296.050 4.280 ;
        RECT 296.890 4.000 370.110 4.280 ;
        RECT 370.950 4.000 444.170 4.280 ;
        RECT 445.010 4.000 518.230 4.280 ;
        RECT 519.070 4.000 592.290 4.280 ;
        RECT 593.130 4.000 647.580 4.280 ;
      LAYER met3 ;
        RECT 4.000 626.640 646.000 643.105 ;
        RECT 4.400 625.240 646.000 626.640 ;
        RECT 4.000 568.840 646.000 625.240 ;
        RECT 4.000 567.440 645.600 568.840 ;
        RECT 4.000 548.440 646.000 567.440 ;
        RECT 4.400 547.040 646.000 548.440 ;
        RECT 4.000 490.640 646.000 547.040 ;
        RECT 4.000 489.240 645.600 490.640 ;
        RECT 4.000 470.240 646.000 489.240 ;
        RECT 4.400 468.840 646.000 470.240 ;
        RECT 4.000 412.440 646.000 468.840 ;
        RECT 4.000 411.040 645.600 412.440 ;
        RECT 4.000 392.040 646.000 411.040 ;
        RECT 4.400 390.640 646.000 392.040 ;
        RECT 4.000 334.240 646.000 390.640 ;
        RECT 4.000 332.840 645.600 334.240 ;
        RECT 4.000 313.840 646.000 332.840 ;
        RECT 4.400 312.440 646.000 313.840 ;
        RECT 4.000 256.040 646.000 312.440 ;
        RECT 4.000 254.640 645.600 256.040 ;
        RECT 4.000 235.640 646.000 254.640 ;
        RECT 4.400 234.240 646.000 235.640 ;
        RECT 4.000 177.840 646.000 234.240 ;
        RECT 4.000 176.440 645.600 177.840 ;
        RECT 4.000 157.440 646.000 176.440 ;
        RECT 4.400 156.040 646.000 157.440 ;
        RECT 4.000 99.640 646.000 156.040 ;
        RECT 4.000 98.240 645.600 99.640 ;
        RECT 4.000 79.240 646.000 98.240 ;
        RECT 4.400 77.840 646.000 79.240 ;
        RECT 4.000 21.440 646.000 77.840 ;
        RECT 4.000 20.040 645.600 21.440 ;
        RECT 4.000 10.715 646.000 20.040 ;
      LAYER met4 ;
        RECT 27.895 637.120 634.505 643.105 ;
        RECT 27.895 117.815 97.440 637.120 ;
        RECT 99.840 117.815 174.240 637.120 ;
        RECT 176.640 117.815 251.040 637.120 ;
        RECT 253.440 117.815 327.840 637.120 ;
        RECT 330.240 117.815 404.640 637.120 ;
        RECT 407.040 117.815 481.440 637.120 ;
        RECT 483.840 117.815 558.240 637.120 ;
        RECT 560.640 117.815 634.505 637.120 ;
  END
END iiitb_rv32i
END LIBRARY

