magic
tech sky130B
magscale 1 2
timestamp 1662902881
<< obsli1 >>
rect 1104 2159 128892 127313
<< obsm1 >>
rect 14 2128 129522 128512
<< metal2 >>
rect 10966 129200 11022 130000
rect 25778 129200 25834 130000
rect 40590 129200 40646 130000
rect 55402 129200 55458 130000
rect 70214 129200 70270 130000
rect 85026 129200 85082 130000
rect 99838 129200 99894 130000
rect 114650 129200 114706 130000
rect 129462 129200 129518 130000
rect 18 0 74 800
rect 14830 0 14886 800
rect 29642 0 29698 800
rect 44454 0 44510 800
rect 59266 0 59322 800
rect 74078 0 74134 800
rect 88890 0 88946 800
rect 103702 0 103758 800
rect 118514 0 118570 800
<< obsm2 >>
rect 20 129144 10910 129200
rect 11078 129144 25722 129200
rect 25890 129144 40534 129200
rect 40702 129144 55346 129200
rect 55514 129144 70158 129200
rect 70326 129144 84970 129200
rect 85138 129144 99782 129200
rect 99950 129144 114594 129200
rect 114762 129144 129406 129200
rect 20 856 129516 129144
rect 130 800 14774 856
rect 14942 800 29586 856
rect 29754 800 44398 856
rect 44566 800 59210 856
rect 59378 800 74022 856
rect 74190 800 88834 856
rect 89002 800 103646 856
rect 103814 800 118458 856
rect 118626 800 129516 856
<< metal3 >>
rect 0 125128 800 125248
rect 129200 113568 130000 113688
rect 0 109488 800 109608
rect 129200 97928 130000 98048
rect 0 93848 800 93968
rect 129200 82288 130000 82408
rect 0 78208 800 78328
rect 129200 66648 130000 66768
rect 0 62568 800 62688
rect 129200 51008 130000 51128
rect 0 46928 800 47048
rect 129200 35368 130000 35488
rect 0 31288 800 31408
rect 129200 19728 130000 19848
rect 0 15648 800 15768
rect 129200 4088 130000 4208
<< obsm3 >>
rect 800 125328 129200 128621
rect 880 125048 129200 125328
rect 800 113768 129200 125048
rect 800 113488 129120 113768
rect 800 109688 129200 113488
rect 880 109408 129200 109688
rect 800 98128 129200 109408
rect 800 97848 129120 98128
rect 800 94048 129200 97848
rect 880 93768 129200 94048
rect 800 82488 129200 93768
rect 800 82208 129120 82488
rect 800 78408 129200 82208
rect 880 78128 129200 78408
rect 800 66848 129200 78128
rect 800 66568 129120 66848
rect 800 62768 129200 66568
rect 880 62488 129200 62768
rect 800 51208 129200 62488
rect 800 50928 129120 51208
rect 800 47128 129200 50928
rect 880 46848 129200 47128
rect 800 35568 129200 46848
rect 800 35288 129120 35568
rect 800 31488 129200 35288
rect 880 31208 129200 31488
rect 800 19928 129200 31208
rect 800 19648 129120 19928
rect 800 15848 129200 19648
rect 880 15568 129200 15848
rect 800 4288 129200 15568
rect 800 4008 129120 4288
rect 800 2143 129200 4008
<< metal4 >>
rect 4208 2128 4528 127344
rect 19568 2128 19888 127344
rect 34928 2128 35248 127344
rect 50288 2128 50608 127344
rect 65648 2128 65968 127344
rect 81008 2128 81328 127344
rect 96368 2128 96688 127344
rect 111728 2128 112048 127344
rect 127088 2128 127408 127344
<< obsm4 >>
rect 5579 127424 126901 128621
rect 5579 23563 19488 127424
rect 19968 23563 34848 127424
rect 35328 23563 50208 127424
rect 50688 23563 65568 127424
rect 66048 23563 80928 127424
rect 81408 23563 96288 127424
rect 96768 23563 111648 127424
rect 112128 23563 126901 127424
<< labels >>
rlabel metal3 s 0 31288 800 31408 6 RN
port 1 nsew signal input
rlabel metal2 s 40590 129200 40646 130000 6 WB_OUT[0]
port 2 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 WB_OUT[10]
port 3 nsew signal output
rlabel metal2 s 114650 129200 114706 130000 6 WB_OUT[11]
port 4 nsew signal output
rlabel metal2 s 10966 129200 11022 130000 6 WB_OUT[12]
port 5 nsew signal output
rlabel metal2 s 99838 129200 99894 130000 6 WB_OUT[13]
port 6 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 WB_OUT[14]
port 7 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 WB_OUT[15]
port 8 nsew signal output
rlabel metal3 s 129200 82288 130000 82408 6 WB_OUT[1]
port 9 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 WB_OUT[2]
port 10 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 WB_OUT[3]
port 11 nsew signal output
rlabel metal3 s 129200 97928 130000 98048 6 WB_OUT[4]
port 12 nsew signal output
rlabel metal3 s 129200 66648 130000 66768 6 WB_OUT[5]
port 13 nsew signal output
rlabel metal2 s 18 0 74 800 6 WB_OUT[6]
port 14 nsew signal output
rlabel metal2 s 85026 129200 85082 130000 6 WB_OUT[7]
port 15 nsew signal output
rlabel metal2 s 25778 129200 25834 130000 6 WB_OUT[8]
port 16 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 WB_OUT[9]
port 17 nsew signal output
rlabel metal3 s 129200 19728 130000 19848 6 clk
port 18 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 io_oeb[0]
port 19 nsew signal output
rlabel metal2 s 129462 129200 129518 130000 6 io_oeb[10]
port 20 nsew signal output
rlabel metal3 s 129200 4088 130000 4208 6 io_oeb[11]
port 21 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 io_oeb[12]
port 22 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_oeb[13]
port 23 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 io_oeb[14]
port 24 nsew signal output
rlabel metal3 s 129200 35368 130000 35488 6 io_oeb[15]
port 25 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 io_oeb[1]
port 26 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 io_oeb[2]
port 27 nsew signal output
rlabel metal3 s 129200 113568 130000 113688 6 io_oeb[3]
port 28 nsew signal output
rlabel metal2 s 55402 129200 55458 130000 6 io_oeb[4]
port 29 nsew signal output
rlabel metal2 s 70214 129200 70270 130000 6 io_oeb[5]
port 30 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 io_oeb[6]
port 31 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 io_oeb[7]
port 32 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 io_oeb[8]
port 33 nsew signal output
rlabel metal3 s 129200 51008 130000 51128 6 io_oeb[9]
port 34 nsew signal output
rlabel metal4 s 4208 2128 4528 127344 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 127344 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 127344 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 127344 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 127344 6 vccd1
port 35 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 127344 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 127344 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 127344 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 127344 6 vssd1
port 36 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 130000 130000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32837506
string GDS_FILE /home/vinay/iiitb_rv32i/openlane/iiitb_rv32i/runs/22_09_11_18_39/results/signoff/iiitb_rv32i.magic.gds
string GDS_START 827710
<< end >>

